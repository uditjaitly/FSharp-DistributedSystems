�      �XMo�8��WpՃm$��=��a�&��"X,�@K��-$7(��w�!��%7N��C��f���������0F+��Q�5\�Q��\9
r��x�0j��9j!�W�G�L��X�,��e���Q����(���l,2�&At�r!����z9ιI�M.�|ِQ �w� �q��*�E��-~K$�G�����7��X%܆s�#n�[Ɠ z�ߎ�X�mD�D��}�|�N%d�s)Yf�#T= ��i�����-S�/�[�z^F<^���y��oU�U��SqWC_�)�<^!E�-!R��)��R젨�WP�|���ӎ΅��?��G�)FjTXa��x9SV�:TƙM? ɐ���2TY��O.�.V���6`@�R����,��[�L��5�dc]��uJ(�G�J�^Xn��=7�����<'D60夙k�f�W��n�TS���k	�,���I�V�>bJ�5!�ck�:�-�.`1@,�i?�ݔ%�(�Bu�ph��y~�KҬS���ڐT/�4��6�iE�ӍDg�/A��36O��{lE�P1��?T��k��ޒ�1%��/7I��OV����؅�p���s�HFx�mj�>���;�~�׺~��p���,pN��\OؔdI�c�:�U�
��Ͻ���*�j롬�w�Ӝ�@k �ũ�@�9�(.���j�?-�J=���\=�T*��HXx+���|M�C:0ޓ�e%�v㴜!�%psFE=��h��B��b�:�_��Z43�o�
�
���+ӄO��q�$z����)��B�@N��N+>?ꍽ�k����қ��j;���{�}�V��r���4��/T�V�>��Jp'C%��V�SC�}t��Y���;D��"��glsB�N`gHS�D�;���S��Wۂu���;�2.�"�V�s��x�F(؊~Rc�bB�/>]|
�d.X��7����;]�2�4KMn&3c.�&0�-�$B>��T2�� ;e�2=��J���/�z,c��q�ZPv���a���S�°��)�x�V|d��b��W��j�D%�3^���ٲm�k�QrzU;����n|9_�(z��q�%[��{G�����t'Į_�/���	�BaP�e���]A4O���>j�&'�K|��
�-���qO�S�����T8I ��dr?�۸�ljBY�mo4�7���H�� �4�����:܋��3�NK,�ݬ�`St��4�9ި#c�O����Y�A�~�}�r��=���L.W)M:`��ަYR7;�����\3�h��P x�2/K�Un�9r=;��^�>�w<�gO�ȼ���i�'�  